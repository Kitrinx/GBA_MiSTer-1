library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity gba_bios is
   port
   (
      clk     : in std_logic;
      address : in std_logic_vector(11 downto 0);
      data    : out std_logic_vector(31 downto 0)
   );
end entity;

architecture arch of gba_bios is

   type t_rom is array(0 to 4095) of std_logic_vector(31 downto 0);
   signal rom : t_rom := ( 
      x"EA000018",
      x"EA000004",
      x"EA00004C",
      x"EA000002",
      x"EA000001",
      x"EA000000",
      x"EA000042",
      x"E59FD1A0",
      x"E92D5000",
      x"E14FC000",
      x"E10FE000",
      x"E92D5000",
      x"E3A0C302",
      x"E5DCE09C",
      x"E35E00A5",
      x"1A000004",
      x"05DCE0B4",
      x"021EE080",
      x"E28FE004",
      x"159FF220",
      x"059FF220",
      x"E59FD164",
      x"E8BD5000",
      x"E169F00C",
      x"E8BD5000",
      x"E25EF004",
      x"E35E0000",
      x"03A0E004",
      x"E3A0C301",
      x"E5DCC300",
      x"E33C0001",
      x"010FC000",
      x"038CC0C0",
      x"0129F00C",
      x"0AFFFFE3",
      x"E3A000DF",
      x"E129F000",
      x"E3A04301",
      x"E5C44208",
      x"EB00000F",
      x"E28F0F96",
      x"E58D00FC",
      x"E59F01CC",
      x"E28FE000",
      x"E12FFF10",
      x"E3A04301",
      x"E5542006",
      x"EB000007",
      x"E3520000",
      x"E9141FFF",
      x"13A0E402",
      x"03A0E302",
      x"E3A0001F",
      x"E129F000",
      x"E3A00000",
      x"E12FFF1E",
      x"E3A000D3",
      x"E129F000",
      x"E59FD0D0",
      x"E3A0E000",
      x"E169F00E",
      x"E3A000D2",
      x"E129F000",
      x"E59FD0B8",
      x"E3A0E000",
      x"E169F00E",
      x"E3A0005F",
      x"E129F000",
      x"E59FD0A0",
      x"E28F0001",
      x"E12FFF10",
      x"49582000",
      x"1D095060",
      x"4770DBFC",
      x"E92D500F",
      x"E3A00301",
      x"E28FE000",
      x"E510F004",
      x"E8BD500F",
      x"E25EF004",
      x"E92D5800",
      x"E55EC002",
      x"E28FB078",
      x"E79BC10C",
      x"E14FB000",
      x"E92D0800",
      x"E20BB080",
      x"E38BB01F",
      x"E129F00B",
      x"E92D4004",
      x"E28FE000",
      x"E12FFF1C",
      x"E8BD4004",
      x"E3A0C0D3",
      x"E129F00C",
      x"E8BD0800",
      x"E169F00B",
      x"E8BD5800",
      x"E1B0F00E",
      x"E3A0C301",
      x"E3A02004",
      x"E5CC2001",
      x"E3A02008",
      x"E5CC2000",
      x"E3A02000",
      x"EA000000",
      x"E3A02080",
      x"E3A0C301",
      x"E5CC2301",
      x"E12FFF1E",
      x"03007F00",
      x"03007FA0",
      x"03007FE0",
      x"03007FF0",
      x"000000B4",
      x"000009C3",
      x"000001A0",
      x"000001A8",
      x"00000330",
      x"00000328",
      x"000003B4",
      x"000003A8",
      x"00000404",
      x"00000474",
      x"000004FD",
      x"00000B4D",
      x"00000BC4",
      x"00000378",
      x"00000C2C",
      x"00000CE0",
      x"00000F60",
      x"000010FC",
      x"00001194",
      x"00001014",
      x"00001279",
      x"000012C1",
      x"00001333",
      x"0000135D",
      x"00001399",
      x"00000801",
      x"00001665",
      x"0000179D",
      x"00001DC5",
      x"0000210D",
      x"00001825",
      x"000018D9",
      x"000013C5",
      x"00001435",
      x"000014C1",
      x"000014FD",
      x"00001515",
      x"000028CF",
      x"0000008C",
      x"000001AC",
      x"00001879",
      x"000018C9",
      x"00002693",
      x"09FE2000",
      x"09FFC000",
      x"00001929",
      x"FFFFFE00",
      x"06242404",
      x"062D2505",
      x"06362606",
      x"20C22100",
      x"32801C22",
      x"72507090",
      x"1C8020FF",
      x"239022A0",
      x"27F09600",
      x"F0009701",
      x"2083FA78",
      x"81A001C0",
      x"62A0480F",
      x"02C01400",
      x"4B0E62E0",
      x"882B602B",
      x"0C624F0D",
      x"80571912",
      x"FA20F003",
      x"70602004",
      x"1BDB7020",
      x"DCF4802B",
      x"900243C8",
      x"A90234D4",
      x"60666021",
      x"60A14901",
      x"FA14F003",
      x"85006000",
      x"FFFFD800",
      x"7FFF7BDE",
      x"00000C63",
      x"E3A03301",
      x"E5932200",
      x"E0022822",
      x"E2121080",
      x"159F07A0",
      x"02021001",
      x"059F079C",
      x"014320B8",
      x"E5C31202",
      x"E12FFF10",
      x"E3A00001",
      x"E3A01001",
      x"E92D4010",
      x"E3A03000",
      x"E3A04001",
      x"E3500000",
      x"1B000004",
      x"E5CC3301",
      x"EB000002",
      x"0AFFFFFC",
      x"E8BD4010",
      x"E12FFF1E",
      x"E3A0C301",
      x"E5CC3208",
      x"E15C20B8",
      x"E0110002",
      x"10222000",
      x"114C20B8",
      x"E5CC4208",
      x"E12FFF1E",
      x"E3A00000",
      x"E3A03000",
      x"E3A0C0DF",
      x"E8B30004",
      x"E129F00C",
      x"E0800002",
      x"E1B01723",
      x"0AFFFFF9",
      x"E12FFF1E",
      x"DC002800",
      x"47704240",
      x"4718A303",
      x"E1A03000",
      x"E1A00001",
      x"E1A01003",
      x"E2113102",
      x"42611000",
      x"E033C040",
      x"22600000",
      x"E1B02001",
      x"E15200A0",
      x"91A02082",
      x"3AFFFFFC",
      x"E1500002",
      x"E0A33003",
      x"20400002",
      x"E1320001",
      x"11A020A2",
      x"1AFFFFF9",
      x"E1A01000",
      x"E1A00003",
      x"E1B0C08C",
      x"22600000",
      x"42611000",
      x"E12FFF1E",
      x"E92D0010",
      x"E1A0C000",
      x"E3A01001",
      x"E1500001",
      x"81A000A0",
      x"81A01081",
      x"8AFFFFFB",
      x"E1A0000C",
      x"E1A04001",
      x"E3A03000",
      x"E1A02001",
      x"E15200A0",
      x"91A02082",
      x"3AFFFFFC",
      x"E1500002",
      x"E0A33003",
      x"20400002",
      x"E1320001",
      x"11A020A2",
      x"1AFFFFF9",
      x"E0811003",
      x"E1B010A1",
      x"E1510004",
      x"3AFFFFEE",
      x"E1A00004",
      x"E8BD0010",
      x"E12FFF1E",
      x"4718A300",
      x"E0010090",
      x"E1A01741",
      x"E2611000",
      x"E3A030A9",
      x"E0030391",
      x"E1A03743",
      x"E2833E39",
      x"E0030391",
      x"E1A03743",
      x"E2833C09",
      x"E283301C",
      x"E0030391",
      x"E1A03743",
      x"E2833C0F",
      x"E28330B6",
      x"E0030391",
      x"E1A03743",
      x"E2833C16",
      x"E28330AA",
      x"E0030391",
      x"E1A03743",
      x"E2833A02",
      x"E2833081",
      x"E0030391",
      x"E1A03743",
      x"E2833C36",
      x"E2833051",
      x"E0030391",
      x"E1A03743",
      x"E2833CA2",
      x"E28330F9",
      x"E0000093",
      x"E1A00840",
      x"E12FFF1E",
      x"2900B5F0",
      x"2800D106",
      x"2000DB01",
      x"2080E049",
      x"E0460200",
      x"D1072800",
      x"DB022900",
      x"02002040",
      x"20C0E03F",
      x"E03C0200",
      x"03921C02",
      x"039B1C0B",
      x"424D4244",
      x"02362640",
      x"29000077",
      x"2800DB1B",
      x"4288DB0F",
      x"1C01DB06",
      x"F7FF1C18",
      x"F7FFFF2D",
      x"E026FF91",
      x"F7FF1C10",
      x"F7FFFF27",
      x"1A30FF8B",
      x"428CE01F",
      x"1C01DBF6",
      x"F7FF1C18",
      x"F7FFFF1D",
      x"1838FF81",
      x"2800E015",
      x"42ACDC09",
      x"1C10DCF3",
      x"FF12F7FF",
      x"FF76F7FF",
      x"1A3019F6",
      x"42A8E009",
      x"1C01DBF5",
      x"F7FF1C18",
      x"F7FFFF07",
      x"19FFFF6B",
      x"BCF01838",
      x"4718BC08",
      x"2608B578",
      x"259E0636",
      x"1E6819AD",
      x"F000211B",
      x"240CF87B",
      x"782B4344",
      x"0F9B079B",
      x"435A2230",
      x"A50918A4",
      x"2400192D",
      x"F0001C20",
      x"2C03F87E",
      x"2C09DB06",
      x"8829DA04",
      x"43310049",
      x"1CAD8808",
      x"2C0B1C64",
      x"BD78D1F0",
      x"7426479B",
      x"6D4F11BC",
      x"32F111BD",
      x"2CE77FD9",
      x"11BD5DA5",
      x"5DA44610",
      x"61734E90",
      x"4E912A84",
      x"75FE106A",
      x"783929C8",
      x"5D1B420E",
      x"12A87838",
      x"67B93F7D",
      x"54EF26F3",
      x"26F27C23",
      x"41376BC6",
      x"730D15AB",
      x"3B4F6BC7",
      x"3DDA5F24",
      x"1749253F",
      x"70E63DDB",
      x"30F7746C",
      x"6738531F",
      x"1A51531E",
      x"5B7D1971",
      x"19704ED6",
      x"75CB3F27",
      x"128C3D62",
      x"2FAD74B8",
      x"64FD74B9",
      x"4F3A6C9A",
      x"73EF276D",
      x"4F3B38B1",
      x"7EA3571E",
      x"35876249",
      x"35861B7C",
      x"67E47AFB",
      x"67E55C92",
      x"438C2BCA",
      x"587F2E6F",
      x"2E6E14B7",
      x"6FA24CB9",
      x"719E38F0",
      x"1F3C475A",
      x"475B6AD8",
      x"32645199",
      x"49EF7B41",
      x"1CD75198",
      x"2403B530",
      x"78022300",
      x"250441E3",
      x"02124053",
      x"DCFB1E6D",
      x"1E491C40",
      x"1C18DCF5",
      x"0F8006C0",
      x"B510BD30",
      x"43442414",
      x"061B2308",
      x"19001D18",
      x"190949F8",
      x"F000220A",
      x"BD10FA33",
      x"49F6B570",
      x"24FF2600",
      x"D1002E98",
      x"2E9A247B",
      x"24FCD100",
      x"DA062E9C",
      x"5D8B5D82",
      x"1C764022",
      x"D0F0429A",
      x"2419E009",
      x"18A45D82",
      x"2EBA1C76",
      x"0620DBFA",
      x"2000D101",
      x"2001E000",
      x"4BE8BD70",
      x"207E2208",
      x"50984240",
      x"2A783210",
      x"4770DBFB",
      x"1EC3B540",
      x"4356009E",
      x"1A9B2340",
      x"1EC0435E",
      x"43432318",
      x"1AF6021B",
      x"2A2F600E",
      x"261ADC07",
      x"3A484356",
      x"23684356",
      x"18F6021B",
      x"BD40604E",
      x"1C0FB5F0",
      x"3680C870",
      x"20801C31",
      x"F7FF0400",
      x"0073FE15",
      x"81FB81BB",
      x"01C9217F",
      x"60796039",
      x"43411221",
      x"31781409",
      x"12298139",
      x"14094341",
      x"81793150",
      x"B5F0BDF0",
      x"9D069C05",
      x"26002700",
      x"184053A0",
      x"42961CB6",
      x"1964DBFA",
      x"429F1C7F",
      x"BDF0DBF5",
      x"2702B5F0",
      x"00434CC2",
      x"19DB181B",
      x"191B009B",
      x"691E685D",
      x"1A5B2320",
      x"434E436B",
      x"095C199B",
      x"0533261F",
      x"0A9D4023",
      x"402302B3",
      x"432B095B",
      x"431C4034",
      x"005E19D3",
      x"18F34BB6",
      x"1E7F801C",
      x"BDF0DAE0",
      x"02092102",
      x"4BB3468C",
      x"4BB2881A",
      x"0D890591",
      x"D0032800",
      x"DA094561",
      x"E0021C92",
      x"DD052900",
      x"801A1E92",
      x"1E522208",
      x"E7E9D5FD",
      x"49AA4770",
      x"01122237",
      x"E00F48A9",
      x"222449A7",
      x"E00B48A8",
      x"06092107",
      x"48A72250",
      x"49A7E006",
      x"D0012800",
      x"18090240",
      x"48A52208",
      x"1852B530",
      x"42984B9B",
      x"2304DB07",
      x"4298031B",
      x"C808DA03",
      x"4291C108",
      x"BD30DBF4",
      x"B085B5F0",
      x"C9A0499D",
      x"C0A0A802",
      x"4B9D489C",
      x"09DB781B",
      x"489CD100",
      x"220A4992",
      x"F95CF000",
      x"FE86F7FF",
      x"1C0B4989",
      x"781833AE",
      x"D0052896",
      x"17D34A96",
      x"A8049304",
      x"F94EF000",
      x"FFBDF7FF",
      x"49934888",
      x"FBAAF000",
      x"49864891",
      x"FC1AF000",
      x"00B82700",
      x"4A839003",
      x"18800238",
      x"02B94B8D",
      x"AA0218C9",
      x"FB40F000",
      x"2F081C7F",
      x"270EDBF1",
      x"4B882403",
      x"19000078",
      x"18C00200",
      x"5BDA4B86",
      x"01214B86",
      x"01891889",
      x"228018C9",
      x"F924F000",
      x"DAEE1E64",
      x"DAEB1EBF",
      x"F000486C",
      x"F000F81C",
      x"F000F82F",
      x"2220F834",
      x"497D9201",
      x"23049100",
      x"497C2204",
      x"F7FF487C",
      x"2105FF38",
      x"43C80609",
      x"20008008",
      x"FF87F7FF",
      x"F7FF2001",
      x"F7FFFF84",
      x"B005FF7D",
      x"B5F1BDF0",
      x"70204C74",
      x"FF72F7FF",
      x"49739800",
      x"F000224E",
      x"485EF8F7",
      x"F0004968",
      x"4867FB55",
      x"60024A6F",
      x"F000495A",
      x"BDF1FD13",
      x"4858B5F1",
      x"4A6C4962",
      x"FAEEF000",
      x"B5F1BDF1",
      x"4C6A4E5F",
      x"25342702",
      x"C40FCE0F",
      x"DCFB1E6D",
      x"1E7F34C0",
      x"2703DCF7",
      x"486502BB",
      x"496518C0",
      x"220118C9",
      x"F0000212",
      x"1E7FF909",
      x"4668DCF4",
      x"49486007",
      x"02122208",
      x"F879F000",
      x"B5F0BDF1",
      x"1C07B081",
      x"24044D5C",
      x"23000624",
      x"21809300",
      x"26808021",
      x"D01D423E",
      x"19090C61",
      x"F0002208",
      x"3920F863",
      x"804843D0",
      x"19090C21",
      x"1D217408",
      x"F0002208",
      x"1F09F859",
      x"F0002210",
      x"21B0F855",
      x"22181909",
      x"F850F000",
      x"0CA0620A",
      x"86208420",
      x"86E084E0",
      x"49492620",
      x"F0002208",
      x"0AE2F845",
      x"3110808A",
      x"700A2207",
      x"F83EF000",
      x"423E2640",
      x"2180D019",
      x"48421909",
      x"71097108",
      x"89086008",
      x"0D800580",
      x"39108108",
      x"31207009",
      x"F0002208",
      x"3940F82B",
      x"3120700A",
      x"F0002208",
      x"2200F825",
      x"19092180",
      x"2601710A",
      x"0AA20861",
      x"F81CF000",
      x"21062608",
      x"0B0A0609",
      x"F816F000",
      x"21072610",
      x"0CA20609",
      x"F810F000",
      x"21052604",
      x"0CA20609",
      x"F80AF000",
      x"21032602",
      x"4A2A0609",
      x"F804F000",
      x"BCF0B001",
      x"4718BC08",
      x"D100423E",
      x"46684770",
      x"E083432A",
      x"00002D71",
      x"0000210D",
      x"03000088",
      x"00003290",
      x"03003580",
      x"00003200",
      x"05000200",
      x"04000088",
      x"03000564",
      x"0000332C",
      x"0000326C",
      x"0000369C",
      x"05000038",
      x"00003264",
      x"000030C0",
      x"0BFE1FE0",
      x"080000B4",
      x"0BFFFFE0",
      x"85000027",
      x"03001564",
      x"06000040",
      x"000030B0",
      x"06010000",
      x"0600B880",
      x"00000202",
      x"00007271",
      x"03007FF7",
      x"03000588",
      x"0000D082",
      x"000030C8",
      x"060024C0",
      x"06002040",
      x"06016800",
      x"85000000",
      x"04000110",
      x"880E0000",
      x"00001F80",
      x"02D4B530",
      x"F0000A64",
      x"D01EF823",
      x"0ED32500",
      x"190DD30C",
      x"D3040E53",
      x"42A9C808",
      x"C108DA15",
      x"42A9E7FB",
      x"C808DA11",
      x"E7FAC108",
      x"0E530864",
      x"8803D305",
      x"DA0842A5",
      x"1CAD534B",
      x"42A5E7FA",
      x"5B43DA03",
      x"1CAD534B",
      x"BC30E7F9",
      x"4718BC08",
      x"46A4A301",
      x"00004718",
      x"E35C0000",
      x"0A000003",
      x"E3CCC4FE",
      x"E080C00C",
      x"E310040E",
      x"131C040E",
      x"E12FFF1E",
      x"4718467B",
      x"E92D47F0",
      x"E1A0A582",
      x"E1B0C4AA",
      x"EBFFFFF3",
      x"0A000012",
      x"E081A4AA",
      x"E1B02CA2",
      x"3A00000B",
      x"E5902000",
      x"E1A03002",
      x"E1A04002",
      x"E1A05002",
      x"E1A06002",
      x"E1A07002",
      x"E1A08002",
      x"E1A09002",
      x"E151000A",
      x"B8A103FC",
      x"BAFFFFFC",
      x"EA000003",
      x"E151000A",
      x"B8B003FC",
      x"B8A103FC",
      x"BAFFFFFB",
      x"E8BD47F0",
      x"E12FFF1E",
      x"E92D0FF0",
      x"E2522001",
      x"BA000027",
      x"E1D031B0",
      x"E1A03423",
      x"E28FCF45",
      x"E2838040",
      x"E20880FF",
      x"E1A08088",
      x"E198B0FC",
      x"E1A08083",
      x"E198C0FC",
      x"E1D090FC",
      x"E1D0A0FE",
      x"E008099B",
      x"E1A03748",
      x"E008099C",
      x"E1A04748",
      x"E0080A9C",
      x"E1A05748",
      x"E0080A9B",
      x"E1A06748",
      x"E8901600",
      x"E1A0B80C",
      x"E1A0B84B",
      x"E1A0C84C",
      x"E26B8000",
      x"E0299893",
      x"E0289C94",
      x"E5818008",
      x"E26B8000",
      x"E02AA895",
      x"E26C8000",
      x"E028A896",
      x"E581800C",
      x"E1C130B0",
      x"E2644000",
      x"E1C140B2",
      x"E1C150B4",
      x"E1C160B6",
      x"E2800014",
      x"E2811010",
      x"EAFFFFD5",
      x"E8BD0FF0",
      x"E12FFF1E",
      x"E92D0F00",
      x"E2522001",
      x"BA000019",
      x"E1D090B4",
      x"E1A09429",
      x"E28FC060",
      x"E2898040",
      x"E20880FF",
      x"E1A08088",
      x"E198B0FC",
      x"E1A08089",
      x"E198C0FC",
      x"E1D090F0",
      x"E1D0A0F2",
      x"E008099B",
      x"E1A08748",
      x"E08180B3",
      x"E008099C",
      x"E1A08748",
      x"E2688000",
      x"E08180B3",
      x"E0080A9C",
      x"E1A08748",
      x"E08180B3",
      x"E0080A9B",
      x"E1A08748",
      x"E08180B3",
      x"E2800008",
      x"EAFFFFE3",
      x"E8BD0F00",
      x"E12FFF1E",
      x"01920000",
      x"04B50323",
      x"07D50645",
      x"0AF10964",
      x"0E050C7C",
      x"11110F8C",
      x"14131294",
      x"1708158F",
      x"19EF187D",
      x"1CC61B5D",
      x"1F8B1E2B",
      x"223D20E7",
      x"24DA238E",
      x"275F261F",
      x"29CD2899",
      x"2C212AFA",
      x"2E5A2D41",
      x"30762F6B",
      x"32743179",
      x"34533367",
      x"36123536",
      x"37AF36E5",
      x"392A3871",
      x"3A8239DA",
      x"3BB63B20",
      x"3CC53C42",
      x"3DAE3D3E",
      x"3E713E14",
      x"3F0E3EC5",
      x"3F843F4E",
      x"3FD33FB1",
      x"3FFB3FEC",
      x"3FFB4000",
      x"3FD33FEC",
      x"3F843FB1",
      x"3F0E3F4E",
      x"3E713EC5",
      x"3DAE3E14",
      x"3CC53D3E",
      x"3BB63C42",
      x"3A823B20",
      x"392A39DA",
      x"37AF3871",
      x"361236E5",
      x"34533536",
      x"32743367",
      x"30763179",
      x"2E5A2F6B",
      x"2C212D41",
      x"29CD2AFA",
      x"275F2899",
      x"24DA261F",
      x"223D238E",
      x"1F8B20E7",
      x"1CC61E2B",
      x"19EF1B5D",
      x"1708187D",
      x"1413158F",
      x"11111294",
      x"0E050F8C",
      x"0AF10C7C",
      x"07D50964",
      x"04B50645",
      x"01920323",
      x"FE6E0000",
      x"FB4BFCDD",
      x"F82BF9BB",
      x"F50FF69C",
      x"F1FBF384",
      x"EEEFF074",
      x"EBEDED6C",
      x"E8F8EA71",
      x"E611E783",
      x"E33AE4A3",
      x"E075E1D5",
      x"DDC3DF19",
      x"DB26DC72",
      x"D8A1D9E1",
      x"D633D767",
      x"D3DFD506",
      x"D1A6D2BF",
      x"CF8AD095",
      x"CD8CCE87",
      x"CBADCC99",
      x"C9EECACA",
      x"C851C91B",
      x"C6D6C78F",
      x"C57EC626",
      x"C44AC4E0",
      x"C33BC3BE",
      x"C252C2C2",
      x"C18FC1EC",
      x"C0F2C13B",
      x"C07CC0B2",
      x"C02DC04F",
      x"C005C014",
      x"C005C000",
      x"C02DC014",
      x"C07CC04F",
      x"C0F2C0B2",
      x"C18FC13B",
      x"C252C1EC",
      x"C33BC2C2",
      x"C44AC3BE",
      x"C57EC4E0",
      x"C6D6C626",
      x"C851C78F",
      x"C9EEC91B",
      x"CBADCACA",
      x"CD8CCC99",
      x"CF8ACE87",
      x"D1A6D095",
      x"D3DFD2BF",
      x"D633D506",
      x"D8A1D767",
      x"DB26D9E1",
      x"DDC3DC72",
      x"E075DF19",
      x"E33AE1D5",
      x"E611E4A3",
      x"E8F8E783",
      x"EBEDEA71",
      x"EEEFED6C",
      x"F1FBF074",
      x"F50FF384",
      x"F82BF69C",
      x"FB4BF9BB",
      x"FE6EFCDD",
      x"4718467B",
      x"E92D4FF0",
      x"E24DD008",
      x"E1D270B0",
      x"E1B0C007",
      x"EBFFFF0B",
      x"0A000022",
      x"E5D26002",
      x"E266A008",
      x"E3A0E000",
      x"E592B004",
      x"E1A08FAB",
      x"E592B004",
      x"E1A0B08B",
      x"E1A0B0AB",
      x"E58DB004",
      x"E5D22003",
      x"E3A03000",
      x"E2577001",
      x"BA000015",
      x"E3A0B0FF",
      x"E1A05A5B",
      x"E4D09001",
      x"E3A04000",
      x"E3540008",
      x"AAFFFFF7",
      x"E009B005",
      x"E1B0C43B",
      x"03580000",
      x"0A000001",
      x"E59DB004",
      x"E08CC00B",
      x"E18EE31C",
      x"E0833002",
      x"E3530020",
      x"BA000002",
      x"E481E004",
      x"E3A0E000",
      x"E3A03000",
      x"E1A05615",
      x"E0844006",
      x"EAFFFFED",
      x"E28DD008",
      x"E8BD4FF0",
      x"E12FFF1E",
      x"4718467B",
      x"E92D4FF0",
      x"E24DD008",
      x"E3B0C402",
      x"EBFFFEDF",
      x"0A000030",
      x"E2802004",
      x"E2827001",
      x"E5D0A000",
      x"E20A400F",
      x"E3A03000",
      x"E3A0E000",
      x"E204A007",
      x"E28AB004",
      x"E58DB004",
      x"E590A000",
      x"E1A0C42A",
      x"E5D2A000",
      x"E28AA001",
      x"E082008A",
      x"E1A02007",
      x"E35C0000",
      x"DA00001F",
      x"E3A08020",
      x"E4905004",
      x"E2588001",
      x"BAFFFFF9",
      x"E3A0A001",
      x"E00A9FA5",
      x"E5D26000",
      x"E1A06916",
      x"E1A0A0A2",
      x"E1A0A08A",
      x"E5D2B000",
      x"E20BB03F",
      x"E28BB001",
      x"E08AA08B",
      x"E08A2009",
      x"E3160080",
      x"0A00000A",
      x"E1A03433",
      x"E5D2A000",
      x"E264B020",
      x"E1833B1A",
      x"E1A02007",
      x"E28EE001",
      x"E59DB004",
      x"E15E000B",
      x"04813004",
      x"024CC004",
      x"03A0E000",
      x"E35C0000",
      x"C1A05085",
      x"CAFFFFE2",
      x"EAFFFFDD",
      x"E28DD008",
      x"E8BD4FF0",
      x"E12FFF1E",
      x"4718467B",
      x"E92D4070",
      x"E4905004",
      x"E1A02425",
      x"E1B0C002",
      x"EBFFFEA4",
      x"0A00001D",
      x"E3520000",
      x"DA00001B",
      x"E4D0E001",
      x"E3A04008",
      x"E2544001",
      x"BAFFFFF9",
      x"E31E0080",
      x"1A000003",
      x"E4D06001",
      x"E4C16001",
      x"E2422001",
      x"EA00000D",
      x"E5D05000",
      x"E3A06003",
      x"E0863245",
      x"E4D06001",
      x"E206500F",
      x"E1A0C405",
      x"E4D06001",
      x"E186500C",
      x"E285C001",
      x"E0422003",
      x"E751500C",
      x"E4C15001",
      x"E2533001",
      x"CAFFFFFB",
      x"E3520000",
      x"C1A0E08E",
      x"CAFFFFE6",
      x"EAFFFFE1",
      x"E8BD4070",
      x"E12FFF1E",
      x"E92D47F0",
      x"E3A03000",
      x"E4908004",
      x"E1A0A428",
      x"E3A02000",
      x"E1B0C00A",
      x"EBFFFE7C",
      x"0A00002E",
      x"E35A0000",
      x"DA00002C",
      x"E4D06001",
      x"E3A07008",
      x"E2577001",
      x"BAFFFFF9",
      x"E3160080",
      x"1A000006",
      x"E4D09001",
      x"E1833219",
      x"E24AA001",
      x"E2322008",
      x"00C130B2",
      x"03A03000",
      x"EA00001B",
      x"E5D09000",
      x"E3A08003",
      x"E0885249",
      x"E4D09001",
      x"E209800F",
      x"E1A04408",
      x"E4D09001",
      x"E1898004",
      x"E2884001",
      x"E2628008",
      x"E2049001",
      x"E028E189",
      x"E04AA005",
      x"E22EE008",
      x"E2628008",
      x"E08481A8",
      x"E1A080A8",
      x"E1A08088",
      x"E11190B8",
      x"E3A080FF",
      x"E0098E18",
      x"E1A08E58",
      x"E1833218",
      x"E2322008",
      x"00C130B2",
      x"03A03000",
      x"E2555001",
      x"CAFFFFF0",
      x"E35A0000",
      x"C1A06086",
      x"CAFFFFD5",
      x"EAFFFFD0",
      x"E8BD47F0",
      x"E12FFF1E",
      x"C808B5F0",
      x"1C3C0A1F",
      x"FC8CF7FF",
      x"2F00D019",
      x"7804DD17",
      x"06621C40",
      x"0A230E52",
      x"1C52D208",
      x"78031ABF",
      x"1C40700B",
      x"1E521C49",
      x"E7EEDCF9",
      x"1ABF1CD2",
      x"1C407805",
      x"1C49700D",
      x"DCFB1E52",
      x"BCF0E7E5",
      x"4718BC08",
      x"B083B5F0",
      x"C8082700",
      x"1C2C0A1D",
      x"FC66F7FF",
      x"2400D02B",
      x"DD282D00",
      x"93017803",
      x"9B011C40",
      x"0E52065A",
      x"0A339E01",
      x"1C52D20E",
      x"78061AAD",
      x"433740A6",
      x"23081C40",
      x"D102405C",
      x"1C89800F",
      x"1E522700",
      x"E7E5DCF3",
      x"1AAD1CD2",
      x"96027806",
      x"9E021C40",
      x"433740A6",
      x"405C2308",
      x"800FD102",
      x"27001C89",
      x"DCF41E52",
      x"B003E7D4",
      x"BC08BCF0",
      x"B5104718",
      x"0A24C810",
      x"FC30F7FF",
      x"7802D00B",
      x"700A1C40",
      x"1E641C49",
      x"7803DD05",
      x"1C40189A",
      x"1C49700A",
      x"BC10E7F7",
      x"4718BC08",
      x"C808B5F0",
      x"1C2C0A1D",
      x"FC1AF7FF",
      x"2408D013",
      x"1C407807",
      x"1E6D1C3A",
      x"7803DD0D",
      x"1C4019DF",
      x"0E36063E",
      x"433240A6",
      x"405C2308",
      x"800AD1F3",
      x"22001C89",
      x"BCF0E7EF",
      x"4718BC08",
      x"C810B510",
      x"F7FF0A24",
      x"D00BFBFD",
      x"1C808802",
      x"1C89800A",
      x"DD051EA4",
      x"189A8803",
      x"800A1C80",
      x"E7F71C89",
      x"BC04BC10",
      x"47084710",
      x"1C14B5B0",
      x"1C071C0D",
      x"DB262A01",
      x"DD002C10",
      x"1C382410",
      x"FFEAF000",
      x"481162FD",
      x"6078723C",
      x"E0042000",
      x"060C1E61",
      x"70280E24",
      x"2C003550",
      x"490CDCF8",
      x"6B094C0C",
      x"42A2680A",
      x"3201D10D",
      x"6A0A600A",
      x"D0032A00",
      x"6A4A63BA",
      x"620863FA",
      x"624F4806",
      x"600C6208",
      x"BCB0637C",
      x"4718BC08",
      x"80000000",
      x"03007FC0",
      x"68736D53",
      x"00002149",
      x"1C07B5F0",
      x"4B206B40",
      x"42981C0C",
      x"3001D138",
      x"21006378",
      x"603C6079",
      x"63386860",
      x"727878A0",
      x"83B82096",
      x"20FF8438",
      x"83F83001",
      x"84B98479",
      x"26006AFD",
      x"1C38E00B",
      x"F0001C29",
      x"20C0FFBA",
      x"00B07028",
      x"68801900",
      x"35506428",
      x"78203601",
      x"DA0B4286",
      x"42B07A38",
      x"E007DCED",
      x"1C291C38",
      x"FFA7F000",
      x"70282000",
      x"36013550",
      x"42B07A38",
      x"78E0DCF4",
      x"D3010A01",
      x"F976F000",
      x"63784802",
      x"BC08BCF0",
      x"00004718",
      x"68736D53",
      x"1C07B5F0",
      x"4E0C6B40",
      x"D11142B0",
      x"63783001",
      x"07F36878",
      x"60784318",
      x"6AFC7A3D",
      x"1C38E005",
      x"F0001C21",
      x"3450FF80",
      x"2D003D01",
      x"637EDCF7",
      x"BC08BCF0",
      x"00004718",
      x"68736D53",
      x"49046B42",
      x"D104428A",
      x"63416842",
      x"08520052",
      x"47706042",
      x"68736D53",
      x"6B47B480",
      x"42974A05",
      x"84C1D105",
      x"21FF8481",
      x"85013101",
      x"BC806342",
      x"00004770",
      x"68736D53",
      x"1C07B5F0",
      x"28008C80",
      x"8CF9D019",
      x"04093901",
      x"84F90C09",
      x"8D39D113",
      x"85393910",
      x"14090409",
      x"DC0F2900",
      x"6AFC7A3D",
      x"E0062600",
      x"1C211C38",
      x"FF3FF000",
      x"34507026",
      x"2D003D01",
      x"BCF0DCF6",
      x"4718BC08",
      x"7A3984F8",
      x"E00A6AF8",
      x"0A137802",
      x"8D3BD305",
      x"74C3089B",
      x"431A2303",
      x"30507002",
      x"29003901",
      x"E7EADCF2",
      x"780DB5B0",
      x"08691C0F",
      x"7CB9D330",
      x"7E3C7CFA",
      x"094A4351",
      x"D1022C01",
      x"56F92316",
      x"2314188A",
      x"004956F9",
      x"56FB2315",
      x"2C0218C9",
      x"2316D102",
      x"185956FB",
      x"42D92380",
      x"4259DA01",
      x"297FE002",
      x"217FDD00",
      x"33791DCB",
      x"0A1B4353",
      x"0E1B061B",
      x"D9002BFF",
      x"743B23FF",
      x"1A59237F",
      x"0A094351",
      x"0E090609",
      x"D90029FF",
      x"747921FF",
      x"D31C08E9",
      x"56F9230E",
      x"43517BFA",
      x"230C0089",
      x"009256FA",
      x"230A1889",
      x"021256FA",
      x"230B1889",
      x"021256FA",
      x"7B7A1889",
      x"7E3A1889",
      x"D1032A00",
      x"56FA2316",
      x"18510112",
      x"723A120A",
      x"4A067279",
      x"6B121C39",
      x"F7FF6BD2",
      x"7838FEB7",
      x"43982305",
      x"BCB07038",
      x"4718BC08",
      x"03007FC0",
      x"1C07B588",
      x"2000491C",
      x"824880C8",
      x"228F481B",
      x"4A1B8082",
      x"7A428042",
      x"0E920692",
      x"431A2340",
      x"011B2335",
      x"18FA7242",
      x"481663C2",
      x"01DB2313",
      x"18F86008",
      x"48146088",
      x"60C84A15",
      x"63074813",
      x"90002000",
      x"1C394668",
      x"FA4EF7FF",
      x"71B82008",
      x"71F8200F",
      x"63B8480F",
      x"62B8480F",
      x"633862F8",
      x"480E63F8",
      x"20016378",
      x"F0000480",
      x"480CF81C",
      x"BC886038",
      x"4718BC08",
      x"040000C0",
      x"04000080",
      x"0000A90E",
      x"040000A0",
      x"040000A4",
      x"03007FC0",
      x"050003EC",
      x"00002425",
      x"00001709",
      x"00003738",
      x"68736D53",
      x"B5904770",
      x"230F491D",
      x"4018041B",
      x"0C006B0F",
      x"491B7238",
      x"18400040",
      x"8BC03820",
      x"01092163",
      x"61381C04",
      x"FFF8F001",
      x"481672F8",
      x"43604B16",
      x"005818C1",
      x"FFF0F001",
      x"06092101",
      x"F0016178",
      x"3001FFEB",
      x"61B81040",
      x"20004C10",
      x"69388060",
      x"F001490F",
      x"2101FFE1",
      x"1A080409",
      x"F0008020",
      x"2001F8AF",
      x"79810680",
      x"D0FC299F",
      x"299F7981",
      x"2080D1FC",
      x"BC908060",
      x"4718BC08",
      x"03007FC0",
      x"000031E8",
      x"00091D1B",
      x"00001388",
      x"04000100",
      x"00044940",
      x"491EB5B0",
      x"6B0F4D1E",
      x"42A96839",
      x"3101D133",
      x"06016039",
      x"D0020E09",
      x"0E490649",
      x"210F7179",
      x"40010209",
      x"0A09D009",
      x"210C71B9",
      x"1DFA2300",
      x"70133249",
      x"39013240",
      x"210FD1FB",
      x"40010309",
      x"0B09D001",
      x"210B71F9",
      x"40010509",
      x"2303D009",
      x"4A0C051B",
      x"7A534019",
      x"069B0B89",
      x"43190E9B",
      x"240F7251",
      x"40040424",
      x"F000D004",
      x"1C20F837",
      x"FF7DF7FF",
      x"BCB0603D",
      x"4718BC08",
      x"03007FC0",
      x"68736D53",
      x"04000080",
      x"4812B5F0",
      x"6B074E12",
      x"42B06838",
      x"3001D11A",
      x"1DF86038",
      x"3049210C",
      x"70022200",
      x"39013040",
      x"DCF92900",
      x"2D0069FD",
      x"2401D00B",
      x"0E000620",
      x"F7FF6AF9",
      x"3401FDB4",
      x"2C043540",
      x"2200DDF6",
      x"603E702A",
      x"BC08BCF0",
      x"00004718",
      x"03007FC0",
      x"68736D53",
      x"480FB588",
      x"6B074B0F",
      x"42986838",
      x"3301D314",
      x"D8114298",
      x"60383001",
      x"490B2000",
      x"80C82335",
      x"71388248",
      x"18F9011B",
      x"46689000",
      x"F7FF4A07",
      x"6838F951",
      x"60383801",
      x"BC08BC88",
      x"00004718",
      x"03007FC0",
      x"68736D53",
      x"040000C0",
      x"05000318",
      x"4802215B",
      x"80C10249",
      x"47708241",
      x"040000C0",
      x"0612B5F0",
      x"29B21C07",
      x"4A0FDD01",
      x"480F21B2",
      x"071C5C43",
      x"00A40F24",
      x"35AD1DC5",
      x"091E592C",
      x"184040F4",
      x"07017840",
      x"00890F09",
      x"09005869",
      x"1B0840C1",
      x"F0001C11",
      x"1901FA51",
      x"F0006878",
      x"BCF0FA4D",
      x"4718BC08",
      x"FF000000",
      x"00003104",
      x"B08DB5F0",
      x"20002100",
      x"20109005",
      x"43CF9003",
      x"910420FF",
      x"F7FF9100",
      x"48FAF840",
      x"70052501",
      x"F7FE2001",
      x"4EF8FF59",
      x"05C12008",
      x"80888035",
      x"0BC088B0",
      x"F7FED001",
      x"F7FEFC91",
      x"20EFFF87",
      x"210101C0",
      x"81C80689",
      x"90022054",
      x"90012076",
      x"02802015",
      x"203B6388",
      x"63C80240",
      x"48EB49EC",
      x"F7FE6108",
      x"F001FECC",
      x"48EAF9EB",
      x"FE66F7FF",
      x"F7FF48E9",
      x"49E9FEFF",
      x"220648E9",
      x"FD0EF7FF",
      x"48E949E8",
      x"F7FF2206",
      x"E156FD09",
      x"E0A82507",
      x"1B422006",
      x"18800090",
      x"42B83008",
      x"DC04920C",
      x"00A94BE2",
      x"3201585A",
      x"4BE0505A",
      x"585A00A9",
      x"01294BDF",
      x"00EC18C9",
      x"92079106",
      x"2307688E",
      x"940B061B",
      x"2E0018E4",
      x"42B8DA67",
      x"3602DC01",
      x"0428608E",
      x"99061400",
      x"FE9AF7FE",
      x"43682014",
      x"184149D4",
      x"9109910A",
      x"F7FE9806",
      x"0168FEA9",
      x"22014BD1",
      x"980918C1",
      x"300C2308",
      x"FE84F001",
      x"42DE2360",
      x"6820DD3E",
      x"430200DA",
      x"43C0203F",
      x"42861C01",
      x"DA016022",
      x"DA1F2D04",
      x"42DE234B",
      x"2E00DB1C",
      x"8820DA13",
      x"03DB2301",
      x"80204318",
      x"4AC2980B",
      x"88A21880",
      x"0A928880",
      x"30040292",
      x"0D800580",
      x"80A04310",
      x"43C0201F",
      x"2303E006",
      x"439A021B",
      x"43C0200F",
      x"60220041",
      x"4BB89A0A",
      x"18108912",
      x"401A6822",
      x"0DC005C0",
      x"43100400",
      x"9A0A6020",
      x"18518952",
      x"02000A00",
      x"0E090609",
      x"60204308",
      x"07014270",
      x"00490F09",
      x"11009A0C",
      x"30010092",
      x"F7FE3201",
      x"9A07FE7D",
      x"38381FD0",
      x"D80C2822",
      x"9A0748A7",
      x"38401880",
      x"68207841",
      x"02120A02",
      x"06001840",
      x"43100E00",
      x"9A076020",
      x"39591FD1",
      x"D80C2950",
      x"F0012005",
      x"3808FE15",
      x"FC50F7FE",
      x"00819A0C",
      x"1C420090",
      x"F7FE2000",
      x"3D01FE59",
      x"E753D400",
      x"06242407",
      x"D0012F6C",
      x"D10D2FB4",
      x"21069802",
      x"90023838",
      x"91049801",
      x"90013880",
      x"9003200A",
      x"4981488F",
      x"E0456108",
      x"DD3F2F6C",
      x"38039802",
      x"98089002",
      x"D1012800",
      x"E0002001",
      x"23032002",
      x"021B6CA1",
      x"07804399",
      x"02000F80",
      x"49824308",
      x"23014001",
      x"18C0049B",
      x"43984B7F",
      x"64A04308",
      x"00E82500",
      x"1DC11900",
      x"22033179",
      x"F7FE1C0E",
      x"8830FFE5",
      x"029B2303",
      x"35014058",
      x"80302D09",
      x"2006DBEF",
      x"F0011C39",
      x"2900FDC3",
      x"9904D109",
      x"31019803",
      x"90033801",
      x"43080200",
      x"49629104",
      x"48708248",
      x"81484960",
      x"E000486F",
      x"2101486F",
      x"80080689",
      x"02009802",
      x"06892101",
      x"98016388",
      x"63C80200",
      x"DB052F10",
      x"F8F4F000",
      x"D1012F10",
      x"E0024967",
      x"D1032FA2",
      x"48574966",
      x"FC22F7FF",
      x"383A1FF8",
      x"D211284F",
      x"28009808",
      x"4862D10E",
      x"6A402301",
      x"D00942D8",
      x"78004860",
      x"D10528F3",
      x"484F495F",
      x"FC0EF7FF",
      x"90082001",
      x"DD0D2F38",
      x"28009808",
      x"9900D00A",
      x"DA022920",
      x"31029900",
      x"221F9100",
      x"99002006",
      x"FDC0F7FE",
      x"FF7AF000",
      x"2001493B",
      x"F0018108",
      x"2F10FD6F",
      x"9904DA09",
      x"31019803",
      x"90033801",
      x"43080200",
      x"49369104",
      x"37018248",
      x"DC002FD2",
      x"484AE6A4",
      x"FD3CF7FE",
      x"1C072600",
      x"4D482800",
      x"9808D102",
      x"D02B2800",
      x"72E82001",
      x"F00071EE",
      x"0600FF55",
      x"72A80E00",
      x"F000D122",
      x"F001F897",
      x"2F00FD47",
      x"79E8D1F3",
      x"D1F02800",
      x"28007AE8",
      x"4838D00B",
      x"43C07800",
      x"401823F3",
      x"4939D0E7",
      x"F7FF4825",
      x"72EEFBBB",
      x"9900E7E1",
      x"DD072900",
      x"221F9900",
      x"91003901",
      x"F7FE2006",
      x"E7D6FD73",
      x"48174931",
      x"61466101",
      x"00CA2100",
      x"230358A7",
      x"439F029B",
      x"29093101",
      x"DBF650A7",
      x"43FF2700",
      x"E00C1C04",
      x"F862F000",
      x"FD12F001",
      x"D2060878",
      x"28109805",
      x"9805D003",
      x"90053001",
      x"37016160",
      x"DDEF2F32",
      x"FDACF7FF",
      x"28007AA8",
      x"20DED03E",
      x"E03BE03D",
      x"04000300",
      x"04000200",
      x"10003F5F",
      x"04000040",
      x"03003B2C",
      x"00940A00",
      x"0300372C",
      x"030036EC",
      x"0300394C",
      x"0300390C",
      x"03003564",
      x"03003580",
      x"030035F0",
      x"07000026",
      x"0000369C",
      x"FE00FFFF",
      x"000036EC",
      x"10001F5F",
      x"00003F27",
      x"00009802",
      x"00001002",
      x"00003908",
      x"000039C0",
      x"03000064",
      x"04000130",
      x"0000389C",
      x"03000088",
      x"03FFFFF0",
      x"00003818",
      x"00103FBF",
      x"F7FE20FF",
      x"B00DFE0C",
      x"BC08BCF0",
      x"00004718",
      x"4710A200",
      x"E0832190",
      x"E2830000",
      x"E12FFF1E",
      x"680048DE",
      x"68034ADE",
      x"D000429A",
      x"1C5B4770",
      x"B5F06003",
      x"464A4641",
      x"465C4653",
      x"B085B41F",
      x"2B006A03",
      x"6A40D003",
      x"F989F000",
      x"6A839805",
      x"F985F000",
      x"69039805",
      x"4DC14698",
      x"7904182D",
      x"D9041E67",
      x"1BC97AC1",
      x"434A4642",
      x"950218AD",
      x"79434EBC",
      x"D02B2B00",
      x"4708A100",
      x"E3540002",
      x"02807E35",
      x"10857008",
      x"E1A04008",
      x"E19500D6",
      x"E1D510D0",
      x"E0800001",
      x"E19710D6",
      x"E0800001",
      x"E0D710D1",
      x"E0800001",
      x"E0010390",
      x"E1A004C1",
      x"E3100080",
      x"12800001",
      x"E7C50006",
      x"E4C50001",
      x"E2544001",
      x"CAFFFFF0",
      x"E28F002F",
      x"E12FFF10",
      x"46412000",
      x"08C91976",
      x"C501D301",
      x"0849C601",
      x"C501D303",
      x"C501C601",
      x"C501C601",
      x"C501C601",
      x"C501C601",
      x"C501C601",
      x"1E49C601",
      x"9C05DCF5",
      x"46816960",
      x"468469A0",
      x"345079A0",
      x"6A639001",
      x"20C77826",
      x"D1004230",
      x"2080E112",
      x"D0144230",
      x"42302040",
      x"2603D119",
      x"1C187026",
      x"62A03010",
      x"61A068D8",
      x"72652500",
      x"78DA61E5",
      x"421020C0",
      x"2010D02F",
      x"70264306",
      x"7A65E02B",
      x"42302004",
      x"7B60D006",
      x"73601E40",
      x"2000D82A",
      x"E0EF7020",
      x"42302040",
      x"79E0D00C",
      x"0A2D4345",
      x"42857B20",
      x"7B25D81E",
      x"D0F02D00",
      x"43062004",
      x"E0177026",
      x"40322203",
      x"D10A2A02",
      x"43457960",
      x"79A00A2D",
      x"D80D4285",
      x"D0EC1C05",
      x"70261E76",
      x"2A03E008",
      x"7920D106",
      x"2DFF182D",
      x"25FFD302",
      x"70261E76",
      x"98057265",
      x"1C4079C0",
      x"09054368",
      x"436878A0",
      x"72A00A00",
      x"436878E0",
      x"72E00A00",
      x"40302010",
      x"D0079004",
      x"30101C18",
      x"18406899",
      x"68D89003",
      x"90041A40",
      x"69A29D02",
      x"A0016AA3",
      x"00004700",
      x"E58D8000",
      x"E5D4A00A",
      x"E5D4B00B",
      x"E5D40001",
      x"E3100008",
      x"0A000013",
      x"E0D360D1",
      x"E0010B96",
      x"E5D50630",
      x"E0800441",
      x"E5C50630",
      x"E0010A96",
      x"E5D50000",
      x"E0800441",
      x"E4C50001",
      x"E2522001",
      x"1A000005",
      x"E59D2010",
      x"E3520000",
      x"159D300C",
      x"1A000001",
      x"E5C42000",
      x"EA000039",
      x"E2588001",
      x"CAFFFFEC",
      x"EA000034",
      x"E594701C",
      x"E594E020",
      x"E1570109",
      x"3A000006",
      x"E3520004",
      x"DA00000D",
      x"E2422004",
      x"E2833004",
      x"E0477109",
      x"E1570109",
      x"2AFFFFF8",
      x"E1570089",
      x"3A000004",
      x"E3520002",
      x"DA000004",
      x"E2422002",
      x"E2833002",
      x"E0477089",
      x"E1570009",
      x"3A00000B",
      x"E2522001",
      x"1A000005",
      x"E59D2010",
      x"E3520000",
      x"159D300C",
      x"1A000002",
      x"E5C42000",
      x"EA00001A",
      x"E2833001",
      x"E0477009",
      x"E1570009",
      x"2AFFFFF3",
      x"E1D300D0",
      x"E1D310D1",
      x"E0411000",
      x"E0060791",
      x"E0010C96",
      x"E0806BC1",
      x"E0010B96",
      x"E5D50630",
      x"E0800441",
      x"E5C50630",
      x"E0010A96",
      x"E5D50000",
      x"E0800441",
      x"E4C50001",
      x"E087700E",
      x"E2588001",
      x"0A000002",
      x"E1570009",
      x"3AFFFFEC",
      x"EAFFFFCD",
      x"E584701C",
      x"E5842018",
      x"E5843028",
      x"E59D8000",
      x"E28F0001",
      x"E12FFF10",
      x"1E409801",
      x"3440DD01",
      x"9805E6E0",
      x"60034B14",
      x"BCFFB006",
      x"46894680",
      x"469B4692",
      x"4718BC08",
      x"00000350",
      x"00000630",
      x"6800480C",
      x"68034A0C",
      x"D10E429A",
      x"1E497901",
      x"DC0A7101",
      x"71017AC1",
      x"21B62000",
      x"4A030209",
      x"80104B03",
      x"80118018",
      x"47708019",
      x"040000C6",
      x"040000D2",
      x"03007FF0",
      x"68736D53",
      x"6B434A98",
      x"D000429A",
      x"1C5B4770",
      x"B5F06343",
      x"464D4644",
      x"465F4656",
      x"1C07B4F0",
      x"2B006BBB",
      x"6BF8D002",
      x"FFC9F7FF",
      x"28006878",
      x"E10CDA00",
      x"6800488B",
      x"1C384680",
      x"F9D8F7FF",
      x"8C398C78",
      x"E0A41840",
      x"6AFD7A3A",
      x"24002301",
      x"21807828",
      x"D1004201",
      x"4691E08B",
      x"431C469A",
      x"6A2C46A3",
      x"D0132C00",
      x"20C77821",
      x"D0094208",
      x"28007C20",
      x"1E40D009",
      x"D1067420",
      x"43012040",
      x"E0027021",
      x"F0001C20",
      x"6B64F8FC",
      x"D1EB2C00",
      x"2040782B",
      x"D03B4218",
      x"F0001C28",
      x"2080F8E7",
      x"20027028",
      x"204073E8",
      x"201674E8",
      x"20017668",
      x"77881DA9",
      x"6C2AE02C",
      x"29807811",
      x"79E9D201",
      x"1C52E004",
      x"29BD642A",
      x"71E9D300",
      x"D30829CF",
      x"6B834640",
      x"38CF1C08",
      x"1C2A1C39",
      x"FF6FF7FF",
      x"29B0E016",
      x"1C08D90F",
      x"72B838B1",
      x"6B5B4643",
      x"181B0080",
      x"1C38681B",
      x"F7FF1C29",
      x"7828FF60",
      x"D0332800",
      x"4856E004",
      x"18093980",
      x"70687808",
      x"28007868",
      x"1E40D0CF",
      x"7E697068",
      x"D0252900",
      x"28007DE8",
      x"7F28D022",
      x"D0022800",
      x"77281E40",
      x"7EA8E01C",
      x"76A81840",
      x"38401C01",
      x"D5020600",
      x"1612060A",
      x"2080E001",
      x"7DE81A42",
      x"11824350",
      x"40507DA8",
      x"D0090600",
      x"782875AA",
      x"29007E29",
      x"210CD101",
      x"2103E000",
      x"70284308",
      x"4653464A",
      x"1E52465C",
      x"2050DD03",
      x"005B182D",
      x"465EE768",
      x"D1032E00",
      x"06002080",
      x"E0606078",
      x"8C78607E",
      x"84783896",
      x"D3002896",
      x"7A3AE756",
      x"78286AFD",
      x"42012180",
      x"210FD04E",
      x"D04B4201",
      x"1C384691",
      x"F7FF1C29",
      x"6A2CF951",
      x"D03E2C00",
      x"20C77821",
      x"D1034208",
      x"F0001C20",
      x"E033F85C",
      x"26077860",
      x"782B4006",
      x"42182003",
      x"7CA1D00E",
      x"43487C28",
      x"70A011C0",
      x"43487C68",
      x"70E011C0",
      x"D0032E00",
      x"21017F60",
      x"77604308",
      x"4218200C",
      x"7A21D01A",
      x"56282008",
      x"D500180A",
      x"2E002200",
      x"4640D00C",
      x"1C116B03",
      x"1C307A6A",
      x"FED1F7FF",
      x"7F606220",
      x"43082102",
      x"E0057760",
      x"7A6A1C11",
      x"F7FF6A60",
      x"6220FAB1",
      x"2C006B64",
      x"7828D1C0",
      x"400821F0",
      x"464A7028",
      x"DD021E52",
      x"182D2050",
      x"4806DCA7",
      x"BCFF6378",
      x"46894680",
      x"469B4692",
      x"4700BC01",
      x"000030D0",
      x"03007FF0",
      x"68736D53",
      x"210046A4",
      x"23002200",
      x"C01E2400",
      x"C01EC01E",
      x"4664C01E",
      x"6AC34770",
      x"D00B2B00",
      x"6B026B41",
      x"D0012A00",
      x"E0006351",
      x"29006219",
      x"630AD000",
      x"62C12100",
      x"B5704770",
      x"78291C0D",
      x"42082080",
      x"6A2CD015",
      x"D0112C00",
      x"78202600",
      x"D00A2800",
      x"23077860",
      x"D0044018",
      x"681B4B85",
      x"F7FF6ADB",
      x"7026FE78",
      x"6B6462E6",
      x"D1EE2C00",
      x"BC70622C",
      x"4700BC01",
      x"4644B5F0",
      x"4656464D",
      x"B4F0465F",
      x"9100B085",
      x"497A1C15",
      x"91016809",
      x"18404979",
      x"71287800",
      x"78186C2B",
      x"D20E2880",
      x"1C5B7168",
      x"28807818",
      x"71A8D208",
      x"78181C5B",
      x"D2032880",
      x"18097929",
      x"1C5B7129",
      x"1C2C642B",
      x"78223424",
      x"421020C0",
      x"796BD024",
      x"42102040",
      x"6AE9D003",
      x"780818C9",
      x"1C18E000",
      x"18090041",
      x"6AA80089",
      x"46891809",
      x"7831464E",
      x"420820C0",
      x"E0B6D000",
      x"42102080",
      x"78F1D00E",
      x"42082080",
      x"39C0D006",
      x"75690049",
      x"21037828",
      x"70284308",
      x"E0017873",
      x"796B46A1",
      x"9E009302",
      x"7F687A71",
      x"28FF1840",
      x"20FFD900",
      x"464E9004",
      x"26077830",
      x"96034006",
      x"9801D018",
      x"2C0069C4",
      x"E090D100",
      x"01B01E76",
      x"78211824",
      x"420820C7",
      x"2040D036",
      x"D1334208",
      x"98047CE1",
      x"D32F4281",
      x"E080D000",
      x"42A86AE0",
      x"E07CD22A",
      x"1C2F9E04",
      x"46902200",
      x"79A39C01",
      x"78213450",
      x"420820C7",
      x"2040D01E",
      x"D0054208",
      x"D1052A00",
      x"7CE61C52",
      x"E00E6AE7",
      x"D10D2A00",
      x"42B07CE0",
      x"1C06D202",
      x"E0066AE7",
      x"6AE0D806",
      x"D90142B8",
      x"E0001C07",
      x"46A0D300",
      x"1E5B3440",
      x"4644DCDF",
      x"D0522C00",
      x"F7FF1C20",
      x"2100FF2C",
      x"6A2B6321",
      x"2B006363",
      x"631CD000",
      x"62E5622C",
      x"77287EE8",
      x"D0014288",
      x"75A976A9",
      x"1C299800",
      x"F804F7FF",
      x"61206868",
      x"74E09804",
      x"72209802",
      x"7830464E",
      x"68777060",
      x"68B06267",
      x"8BE86060",
      x"7CA181A0",
      x"43487C28",
      x"70A011C0",
      x"43487C68",
      x"70E011C0",
      x"20087A21",
      x"180B5628",
      x"2300D500",
      x"2E009E03",
      x"464ED00F",
      x"77A078B0",
      x"208078F1",
      x"D1004208",
      x"7A6A77E1",
      x"98031C19",
      x"6B1B9B01",
      x"FD87F7FF",
      x"7A6AE004",
      x"1C381C19",
      x"F96CF7FF",
      x"20806220",
      x"78297020",
      x"400820F0",
      x"B0057028",
      x"4680BCFF",
      x"46924689",
      x"BC01469B",
      x"00004700",
      x"03007FF0",
      x"000030D0",
      x"6C0AB510",
      x"2B807813",
      x"714BD203",
      x"640A1C52",
      x"794BE000",
      x"29006A09",
      x"2483D00D",
      x"4222780A",
      x"7C48D006",
      x"D1034298",
      x"43022040",
      x"E002700A",
      x"29006B49",
      x"BC10D1F2",
      x"4700BC01",
      x"1C0DB530",
      x"2C006A2C",
      x"7821D00C",
      x"420820C7",
      x"2040D002",
      x"70214301",
      x"F7FF1C20",
      x"6B64FEA2",
      x"D1F22C00",
      x"70282000",
      x"BC01BC30",
      x"46F44700",
      x"4A0A2124",
      x"F0006813",
      x"C008F806",
      x"1E491D12",
      x"4760DCF8",
      x"B4017813",
      x"D1050E50",
      x"42824803",
      x"0B90D301",
      x"2300D000",
      x"4770BC01",
      x"00003738",
      x"1C536C0A",
      x"7813640B",
      x"B500E7ED",
      x"78D06C0A",
      x"78930200",
      x"02004318",
      x"43187853",
      x"F7FF0200",
      x"4318FFE1",
      x"BC016408",
      x"788A4700",
      x"D2082A03",
      x"188B0092",
      x"1D126C0A",
      x"788A645A",
      x"708A1C52",
      x"E7ADE7E3",
      x"2A00788A",
      x"1E52D005",
      x"0092708A",
      x"6C5A188B",
      x"4770640A",
      x"6C0AB500",
      x"2B007813",
      x"1C52D102",
      x"E7D1640A",
      x"1C5B78CB",
      x"469C70CB",
      x"FFC6F7FF",
      x"D200459C",
      x"2300E7C8",
      x"1D5270CB",
      x"BC01640A",
      x"46F44700",
      x"FFBAF7FF",
      x"4760774B",
      x"F7FF46F4",
      x"005BFFB5",
      x"8BC28383",
      x"0A1B4353",
      x"47608403",
      x"F7FF46F4",
      x"728BFFAB",
      x"220C780B",
      x"700B4313",
      x"46F44760",
      x"78136C0A",
      x"640A1C52",
      x"18D2005A",
      x"6B030092",
      x"681318D2",
      x"FF8BF7FF",
      x"6853624B",
      x"FF87F7FF",
      x"6893628B",
      x"FF83F7FF",
      x"476062CB",
      x"F7FF46F4",
      x"748BFF8B",
      x"2203780B",
      x"700B4313",
      x"46F44760",
      x"FF82F7FF",
      x"750B3B40",
      x"2203780B",
      x"700B4313",
      x"46F44760",
      x"FF78F7FF",
      x"738B3B40",
      x"220C780B",
      x"700B4313",
      x"46F44760",
      x"FF6EF7FF",
      x"780B73CB",
      x"4313220C",
      x"4760700B",
      x"F7FF46F4",
      x"764BFF65",
      x"D1002B00",
      x"4760758B",
      x"F7FF46F4",
      x"76CBFF5D",
      x"46F44760",
      x"FF58F7FF",
      x"2B0075CB",
      x"758BD100",
      x"46F44760",
      x"FF50F7FF",
      x"42987E08",
      x"760BD004",
      x"220F780B",
      x"700B4313",
      x"46F44760",
      x"FF44F7FF",
      x"730B3B40",
      x"220C780B",
      x"700B4313",
      x"46F44760",
      x"78136C0A",
      x"48031C52",
      x"F7FF18C0",
      x"7003FF36",
      x"00004760",
      x"04000060",
      x"1C292620",
      x"086D4051",
      x"D3000849",
      x"08524045",
      x"D1F61E76",
      x"B5544770",
      x"657B468C",
      x"6BB96C7B",
      x"10891AC9",
      x"2989DD17",
      x"2189DD00",
      x"8C3D687C",
      x"46616539",
      x"1C64434C",
      x"4062681A",
      x"404A4259",
      x"404A6D79",
      x"847DC304",
      x"FFDAF7FF",
      x"1E496D39",
      x"843DD1EE",
      x"BD54607C",
      x"F000B500",
      x"BC02F8F2",
      x"8931468E",
      x"D2FC0A09",
      x"B5FA4770",
      x"A2CB23DF",
      x"F8E6F000",
      x"24FF1C07",
      x"F95EF7FE",
      x"0D3CD045",
      x"402323E8",
      x"D1402B20",
      x"29012400",
      x"2902D003",
      x"4CC8DC3B",
      x"877C430C",
      x"61386A38",
      x"1A246A7C",
      x"401C4BC0",
      x"F7FE60FC",
      x"D02EF947",
      x"89604CBE",
      x"43108AE2",
      x"43108C62",
      x"43108DE2",
      x"D2240C00",
      x"7FB84EBA",
      x"0F400700",
      x"8F7A8831",
      x"D0022A00",
      x"0FC007C0",
      x"72387D39",
      x"4BB67139",
      x"49FA0C1B",
      x"4CFB2A00",
      x"49F9D102",
      x"4CFA4BAE",
      x"873B87F9",
      x"69B9643C",
      x"7F396039",
      x"1C347039",
      x"D3050840",
      x"297378E1",
      x"1CA4D101",
      x"E08EE7F8",
      x"68FDD1FB",
      x"383408A8",
      x"19496939",
      x"49A260F9",
      x"D1FD1E49",
      x"FF9AF7FF",
      x"71798871",
      x"88F288B1",
      x"2B008F7B",
      x"21FFD001",
      x"71B922FF",
      x"240271FA",
      x"693B46A4",
      x"1AC96A39",
      x"8FB80889",
      x"681AD217",
      x"8F3D8FF8",
      x"FF56F7FF",
      x"6839873D",
      x"434148E1",
      x"60391C49",
      x"40486818",
      x"1A5A6A39",
      x"185249F1",
      x"6C3A4251",
      x"40484051",
      x"87BA0C02",
      x"F7FF4E8C",
      x"6A39FF72",
      x"D0184299",
      x"1A5C46A6",
      x"8F791EA4",
      x"D0002900",
      x"49E71EA4",
      x"7A3A1864",
      x"08521C35",
      x"8869D305",
      x"04094061",
      x"1CADD141",
      x"D1FCE7F7",
      x"45624674",
      x"2000D101",
      x"F000E03A",
      x"2C00F844",
      x"1C9BD00C",
      x"29008F79",
      x"1C9BD000",
      x"D1022C02",
      x"429968F9",
      x"2065D1B6",
      x"E7D01E64",
      x"F7FF2401",
      x"7A3AFF42",
      x"08521C33",
      x"8859D309",
      x"D0042975",
      x"D11C2865",
      x"D11A2974",
      x"1C9B2400",
      x"D1FCE7F3",
      x"D0052866",
      x"D0002C00",
      x"F0002066",
      x"E7E5F81C",
      x"D00C2C00",
      x"8F3D8FF8",
      x"F7FF687A",
      x"4E64FEF3",
      x"F7FF1C28",
      x"2100FF1B",
      x"1C04468C",
      x"2001E7B5",
      x"63F863B8",
      x"1C396438",
      x"C7013114",
      x"D1FC42B9",
      x"BC04BCFA",
      x"21964710",
      x"D1FD1E49",
      x"81706030",
      x"29008F79",
      x"49B8D100",
      x"47708131",
      x"48B7B500",
      x"29017801",
      x"7AB8D10E",
      x"D30B0640",
      x"7CF97CB8",
      x"D1094308",
      x"49AF6BB8",
      x"DA031A09",
      x"74B82078",
      x"E2A94899",
      x"BD002000",
      x"035168BA",
      x"7D380F89",
      x"1E491CC0",
      x"7538D5FC",
      x"06810880",
      x"40510312",
      x"404817C9",
      x"4001211F",
      x"025068BA",
      x"28070F40",
      x"2100DB05",
      x"0F400310",
      x"DB002807",
      x"221F2000",
      x"FE4CF7FD",
      x"1E407CB8",
      x"74B8DB01",
      x"2005D1DA",
      x"BD0074F8",
      x"B500B4F0",
      x"4C354F99",
      x"49806CF8",
      x"1C404348",
      x"E28064F8",
      x"21E06CF8",
      x"21A04388",
      x"23804048",
      x"4398021B",
      x"780A4990",
      x"D0032A01",
      x"6A4A492E",
      x"D1001C52",
      x"60384318",
      x"7BBE7BFD",
      x"28007B78",
      x"F000D11B",
      x"7B3BF8F1",
      x"2E028A20",
      x"1E5BD104",
      x"2600D510",
      x"E00A2306",
      x"D1042E01",
      x"D5091E5B",
      x"23062602",
      x"1E5BE003",
      x"2601D504",
      x"491C231E",
      x"25006379",
      x"F000733B",
      x"2D00F8DB",
      x"613DD136",
      x"4A6472BD",
      x"4A7663BA",
      x"647A63FA",
      x"73FA2201",
      x"2E0073BE",
      x"22C0D10B",
      x"82A20212",
      x"63656B21",
      x"21078725",
      x"21AD8421",
      x"84390149",
      x"2E01E0B9",
      x"82A5D106",
      x"49074A58",
      x"81658122",
      x"E7F46025",
      x"4ADA82A5",
      x"49070C12",
      x"E7F50C09",
      x"E129F003",
      x"E12FFF1E",
      x"0003FFF8",
      x"040000B0",
      x"04000120",
      x"0000301D",
      x"C3871089",
      x"03000064",
      x"D1192D01",
      x"F89AF000",
      x"80592180",
      x"430A881A",
      x"811D801A",
      x"D1052E00",
      x"84212147",
      x"E007A2C9",
      x"E00349C7",
      x"D1FB2E01",
      x"0C094940",
      x"A2558121",
      x"73F92102",
      x"E07E637A",
      x"D1002D02",
      x"F7FFE07B",
      x"2D03FF2D",
      x"2800D002",
      x"E075D075",
      x"F876F000",
      x"1E406B38",
      x"2E00D509",
      x"8F21D104",
      x"40112230",
      x"E780D004",
      x"D1852E01",
      x"6338E789",
      x"81182001",
      x"28007C78",
      x"2E00D15C",
      x"483FD129",
      x"49F80C00",
      x"F7FF4B26",
      x"647BFDEA",
      x"428B6BF9",
      x"6BB8D153",
      x"D1504058",
      x"880A1F09",
      x"42938C7B",
      x"6008D114",
      x"4AF668B9",
      x"42914011",
      x"7AB9D10E",
      x"18897A3A",
      x"18897A7A",
      x"1A897AFA",
      x"D1050649",
      x"210148F0",
      x"F99DF000",
      x"D0332800",
      x"73F82000",
      x"6BFAE033",
      x"42936C7B",
      x"480ED02F",
      x"2E024B0F",
      x"480BD101",
      x"49104B0C",
      x"FDB9F7FF",
      x"D10C429A",
      x"F7FF69FA",
      x"843DFDA9",
      x"210448E3",
      x"1B897BBE",
      x"F97FF000",
      x"D1E12800",
      x"647B6BFB",
      x"0000E015",
      x"0000C37B",
      x"0000A517",
      x"43202F2F",
      x"6465646F",
      x"20796220",
      x"6177614B",
      x"6F646573",
      x"02000000",
      x"60032003",
      x"74782004",
      x"200073F8",
      x"4718BCF8",
      x"4BCA2000",
      x"47708118",
      x"E7FA2001",
      x"21004BCB",
      x"477073D9",
      x"88114AC1",
      x"7B984BC8",
      x"D1042801",
      x"09C08910",
      x"6B58D26F",
      x"28024687",
      x"8C11D0FB",
      x"20078411",
      x"E7F64001",
      x"020000C0",
      x"A1C12083",
      x"03007FFB",
      x"0300000C",
      x"28620A08",
      x"7B98D16C",
      x"D1012802",
      x"E0022001",
      x"06808910",
      x"75980F80",
      x"2101D051",
      x"75594081",
      x"A00A8811",
      x"74196358",
      x"7318200B",
      x"40082011",
      x"0908D145",
      x"090A4308",
      x"4042404A",
      x"D13E0712",
      x"02002072",
      x"43017D59",
      x"0000E0A7",
      x"28620A08",
      x"2861D0E9",
      x"2003D133",
      x"735873D8",
      x"639A4AA4",
      x"A0012260",
      x"0000E008",
      x"80116B9A",
      x"639A1C92",
      x"1E526C9A",
      x"A003D100",
      x"0212649A",
      x"43117D59",
      x"0000E08A",
      x"28630A08",
      x"20FFD1E1",
      x"76D87698",
      x"76197299",
      x"28027B98",
      x"7DD8D102",
      x"E0057658",
      x"76588850",
      x"76988890",
      x"76D888D0",
      x"60586998",
      x"75DA785A",
      x"2173A002",
      x"43110209",
      x"E078E06C",
      x"28630A08",
      x"2864D0E4",
      x"7719D173",
      x"7B98789A",
      x"D1032802",
      x"20FF775A",
      x"77D87798",
      x"E7EAA001",
      x"0000E05E",
      x"28027B98",
      x"8850D005",
      x"88907758",
      x"88D07798",
      x"008977D8",
      x"487731C8",
      x"40414008",
      x"4979D157",
      x"3208180A",
      x"A00163DA",
      x"0000E044",
      x"28027B98",
      x"80016B98",
      x"6811D102",
      x"1C806001",
      x"63991C81",
      x"42886BD8",
      x"A001D137",
      x"0000E034",
      x"D13E2965",
      x"6BDA6C59",
      x"D0014291",
      x"E02C2174",
      x"A0012175",
      x"0000E028",
      x"D0F92965",
      x"D1302966",
      x"A0018C19",
      x"0000E020",
      x"42888C18",
      x"7B99D129",
      x"D10C2901",
      x"071B7C1B",
      x"085B0F5B",
      x"8851D304",
      x"D1024288",
      x"E7F81C92",
      x"4B5ED1FC",
      x"69D8D119",
      x"1A407E59",
      x"1A407E99",
      x"1A407ED9",
      x"06003811",
      x"21FFD10F",
      x"A0387459",
      x"4A4E6358",
      x"80518151",
      x"28027B98",
      x"4A4BD102",
      x"81104804",
      x"6318200B",
      x"21004770",
      x"A03073D9",
      x"0000E7EE",
      x"10085088",
      x"D1F62901",
      x"60586818",
      x"40484945",
      x"200B6350",
      x"21107318",
      x"E04BA000",
      x"D1EA2904",
      x"73D82003",
      x"A0017358",
      x"0000E046",
      x"D1E22902",
      x"21026B10",
      x"40010209",
      x"A23909C9",
      x"68111852",
      x"60984048",
      x"227F0A01",
      x"04004011",
      x"3180D300",
      x"40100C00",
      x"430101C9",
      x"00C9313F",
      x"4008482F",
      x"D0054288",
      x"06407A98",
      x"72980E40",
      x"01C02089",
      x"4930300C",
      x"64191809",
      x"A0012120",
      x"0000E01A",
      x"D1B82902",
      x"21108F10",
      x"6B104041",
      x"6B998711",
      x"6399C101",
      x"42886BD8",
      x"4924D1A4",
      x"D1024288",
      x"63D86C18",
      x"4822E79E",
      x"68006841",
      x"63504348",
      x"A0022100",
      x"87114A18",
      x"E7936358",
      x"B5004770",
      x"60104A1C",
      x"71194B19",
      x"D0012901",
      x"71587DB8",
      x"F7FD1D10",
      x"BD00FB59",
      x"F7FD1D00",
      x"8CB8FC86",
      x"D1012800",
      x"84B8203C",
      x"7CB8E54E",
      x"D1022877",
      x"FC90F7FD",
      x"2876E003",
      x"F7FDD101",
      x"8CB8FC92",
      x"D0072800",
      x"84B81E40",
      x"D1032839",
      x"490F480E",
      x"F9E0F7FE",
      x"0000E568",
      x"04000120",
      x"0003FFF8",
      x"6177614B",
      x"6F646573",
      x"04000200",
      x"020000C0",
      x"020001F8",
      x"02000000",
      x"0300000C",
      x"80808080",
      x"EA000036",
      x"EA00002E",
      x"0300390C",
      x"00003980",
      x"00280022",
      x"00880082",
      x"00E800E2",
      x"01480142",
      x"08020200",
      x"00000000",
      x"080101C0",
      x"0000001E",
      x"03020100",
      x"07060504",
      x"0B0A0908",
      x"0F0E0D0C",
      x"13121110",
      x"17161514",
      x"201E1C18",
      x"2C2A2824",
      x"38363430",
      x"4442403C",
      x"504E4C48",
      x"5C5A5854",
      x"00000060",
      x"E3E2E1E0",
      x"E7E6E5E4",
      x"EBEAE9E8",
      x"D3D2D1D0",
      x"D7D6D5D4",
      x"DBDAD9D8",
      x"C3C2C1C0",
      x"C7C6C5C4",
      x"CBCAC9C8",
      x"B3B2B1B0",
      x"B7B6B5B4",
      x"BBBAB9B8",
      x"A3A2A1A0",
      x"A7A6A5A4",
      x"ABAAA9A8",
      x"93929190",
      x"97969594",
      x"9B9A9998",
      x"83828180",
      x"87868584",
      x"8B8A8988",
      x"73727170",
      x"77767574",
      x"7B7A7978",
      x"63626160",
      x"67666564",
      x"6B6A6968",
      x"53525150",
      x"57565554",
      x"5B5A5958",
      x"43424140",
      x"47464544",
      x"4B4A4948",
      x"33323130",
      x"37363534",
      x"3B3A3938",
      x"23222120",
      x"27262524",
      x"2B2A2928",
      x"13121110",
      x"17161514",
      x"1B1A1918",
      x"03020100",
      x"07060504",
      x"0B0A0908",
      x"80000000",
      x"879C7C97",
      x"8FACD61E",
      x"9837F052",
      x"A14517CC",
      x"AADC0848",
      x"B504F334",
      x"BFC886BB",
      x"CB2FF52A",
      x"D744FCCB",
      x"E411F03A",
      x"F1A1BF39",
      x"00840060",
      x"00E000B0",
      x"01300108",
      x"01C00160",
      x"02600210",
      x"02C002A0",
      x"FFFFFFFF",
      x"01F0001F",
      x"01F0281F",
      x"01F0581F",
      x"01F00000",
      x"01F0280A",
      x"01F05816",
      x"01F07C00",
      x"01F07C0A",
      x"01F07C16",
      x"00007C00",
      x"00A07C0A",
      x"01607C16",
      x"00007C1F",
      x"00A07C1F",
      x"01607C1F",
      x"0000001F",
      x"00A0281F",
      x"0160581F",
      x"01F0001F",
      x"01F0281F",
      x"01F0581F",
      x"01F07C1F",
      x"01F07C1F",
      x"01F07C1F",
      x"FF1F7C00",
      x"7C1FFD5F",
      x"0000D424",
      x"0000400F",
      x"82810100",
      x"830F8382",
      x"8303C30C",
      x"C3048301",
      x"C2020E08",
      x"0B07C20D",
      x"09050A06",
      x"51AEFF24",
      x"21A29A69",
      x"0A82843D",
      x"AD09E484",
      x"988B2411",
      x"217F81C0",
      x"19BE52A3",
      x"20CE0993",
      x"4A4A4610",
      x"EC3127F8",
      x"33E8C758",
      x"BFCEE382",
      x"94DFF485",
      x"C1094BCE",
      x"C08A5694",
      x"FCA77213",
      x"734D849F",
      x"619ACAA3",
      x"27A39758",
      x"769803FC",
      x"61C71D23",
      x"56AE0403",
      x"008438BF",
      x"FD0EA740",
      x"03FE52FF",
      x"F130956F",
      x"85C0FB97",
      x"2580D660",
      x"03BE63A9",
      x"E2384E01",
      x"FF34A2F9",
      x"44033EBB",
      x"CB900078",
      x"943A1188",
      x"637CC065",
      x"AF3CF087",
      x"8BE425D6",
      x"72AC0A38",
      x"07F8D421",
      x"0003C024",
      x"0180000F",
      x"42014100",
      x"43C20502",
      x"C4430143",
      x"03C30F0A",
      x"09C302C3",
      x"0807040B",
      x"0E0C0D06",
      x"38540300",
      x"481C0C02",
      x"9956C0C3",
      x"756D8008",
      x"441AA6D9",
      x"80844021",
      x"1035B7A6",
      x"F1DB6C98",
      x"66D415A2",
      x"002C0A07",
      x"B1AC0418",
      x"55E19DEB",
      x"45B048DE",
      x"46EC6C1A",
      x"6004D858",
      x"292E0104",
      x"E2AF60C7",
      x"1061D661",
      x"E40FC69D",
      x"40381379",
      x"1B775617",
      x"5AB06E8D",
      x"BC36E230",
      x"C33D6C28",
      x"C1F0E1E7",
      x"B49A9D14",
      x"0AA08094",
      x"56746946",
      x"DA0DB505",
      x"5B043079",
      x"220D1268",
      x"46A51990",
      x"91F0E3D0",
      x"E225724D",
      x"C9401866",
      x"A0AC0618",
      x"83C84C85",
      x"B486F181",
      x"E5D9286D",
      x"6A280AB6",
      x"2F94B1B7",
      x"57A34D5B",
      x"CD1BF87E",
      x"D3AF430D",
      x"FA379A37",
      x"95B69BDA",
      x"B69112C4",
      x"00A85A1D",
      x"79B4A013",
      x"928110D2",
      x"0A86DA46",
      x"88DC30A3",
      x"306CD6C0",
      x"E686F19C",
      x"00C300F4",
      x"161E82C6",
      x"6ABBD060",
      x"24056320",
      x"2BFBA50A",
      x"1B9E5438",
      x"5A909790",
      x"3890DE7F",
      x"0A328283",
      x"8012B5B0",
      x"98C37904",
      x"D03862E3",
      x"DF465D5F",
      x"D91F29C3",
      x"54A1E55F",
      x"CA480069",
      x"6C16ECA3",
      x"B30C3506",
      x"F6ADF5B7",
      x"F0DA065B",
      x"6DBC9BC0",
      x"4B4B69AE",
      x"21870F2A",
      x"100CA45B",
      x"6510AFDA",
      x"5B86DCF2",
      x"B8D11BC3",
      x"E6987A51",
      x"D8B69675",
      x"ADE739DD",
      x"CE37DBE7",
      x"28CFCE74",
      x"5066DCD8",
      x"B6DADB4A",
      x"DBC826A1",
      x"F620D542",
      x"DEE14B19",
      x"AA8D37BA",
      x"BCCCF29C",
      x"B479EEC7",
      x"CF202C02",
      x"D25B4CCE",
      x"8D7ABB63",
      x"0364DAFA",
      x"F999FE70",
      x"7520AA9F",
      x"836F272E",
      x"39F55052",
      x"6EB2587E",
      x"9AF255B9",
      x"8A05DA0D",
      x"BAB079AB",
      x"7EADF5B7",
      x"E8E68F99",
      x"77EE9248",
      x"18851954",
      x"08485CDE",
      x"73685A4C",
      x"8441E67D",
      x"F0D44883",
      x"36BC37B7",
      x"E53A726A",
      x"90999EAE",
      x"2403190A",
      x"F0AE8574",
      x"ECC5AD35",
      x"61BC48DF",
      x"3F4A628F",
      x"93325CCD",
      x"99B3CCAD",
      x"8E650C2A",
      x"BBAA4950",
      x"306D29CB",
      x"5F4E9FA3",
      x"5333746D",
      x"386B15A5",
      x"C62D0996",
      x"8A31F64E",
      x"7EA53DE2",
      x"A8485C24",
      x"31086895",
      x"8B99421C",
      x"18B5C3BB",
      x"9A3BD91C",
      x"CDA2B5DE",
      x"AA776D38",
      x"6F438ED0",
      x"EF4AE4F1",
      x"9C2FA805",
      x"65A50651",
      x"A766EA6C",
      x"FFB3F0D9",
      x"86EE4C37",
      x"B46FAD09",
      x"D069D293",
      x"A4CC2219",
      x"7BBE7CCD",
      x"107CBA0B",
      x"FF2AAB4E",
      x"81079132",
      x"5265A550",
      x"B1733016",
      x"AD046645",
      x"825BAB5A",
      x"ED4884D2",
      x"6429185E",
      x"4BEACB32",
      x"025FBB58",
      x"5AEFDB5C",
      x"AE6D77DA",
      x"4FEBC4DB",
      x"76517466",
      x"156DCB58",
      x"955EF43F",
      x"73A2FA52",
      x"484CE119",
      x"1FCD1934",
      x"D1143998",
      x"77D57FA0",
      x"E51A4A37",
      x"216D2AF6",
      x"A531EC87",
      x"E79F2600",
      x"0502100A",
      x"8108815C",
      x"88222098",
      x"854440B0",
      x"68051581",
      x"D2488844",
      x"5A2442C4",
      x"135AFD91",
      x"1022E832",
      x"22C88044",
      x"88810888",
      x"AC461514",
      x"21AA21C4",
      x"6197C5AA",
      x"64900888",
      x"B4C46B88",
      x"45C4235B",
      x"69882F83",
      x"A59ED758",
      x"8C21159B",
      x"AA70487D",
      x"5A02E967",
      x"B5A62362",
      x"3EC5900D",
      x"421100A8",
      x"0E8298AB",
      x"B9986158",
      x"2FA95019",
      x"4199BEDC",
      x"0B448804",
      x"A1244400",
      x"D45D9088",
      x"74294E00",
      x"00000000",
      x"C2AD2620",
      x"01000A40",
      x"C4962620",
      x"0040098C",
      x"C67F2620",
      x"00000980",
      x"C8682620",
      x"000008CC",
      x"CA502620",
      x"000008C0",
      x"CC392620",
      x"0000080C",
      x"CE222620",
      x"00000800",
      x"C0376466",
      x"00005B40",
      x"C0776466",
      x"00005B50",
      x"81742268",
      x"00000290",
      x"FFFEFEFE",
      x"FF00FFFF",
      x"00010000",
      x"02010101",
      x"FFFF0202",
      x"0000FF00",
      x"01010001",
      x"0000FF00",
      x"00000001",
      x"00004778",
      x"EAFFF2A1",
      x"00004778",
      x"EAFFF29A",
      x"00004778",
      x"EAFFF31F",
      x"00004778",
      x"EAFFF2FD",
      x"00004778",
      x"EAFFF569",
      x"00002665",
      x"000026CF",
      x"000026EF",
      x"00002709",
      x"0000271D",
      x"00002665",
      x"00002665",
      x"00002665",
      x"00002665",
      x"0000274B",
      x"00002755",
      x"00002769",
      x"0000277B",
      x"000027A9",
      x"000027BB",
      x"000027CF",
      x"000027E3",
      x"000027F5",
      x"00002805",
      x"0000280F",
      x"0000281F",
      x"00002665",
      x"00002665",
      x"00002837",
      x"00002665",
      x"00002665",
      x"00002665",
      x"0000284B",
      x"00002665",
      x"00002629",
      x"0000170B",
      x"000023E7",
      x"00001535",
      x"0000159D",
      x"000023C7",
      x"000023B1",
      x"00003C00",
      x"0000382C",
      x"BC4D00FF",
      x"00003C00",
      x"000039D0",
      x"F99AA5FF",
      x"00003C00",
      x"0000382C",
      x"F680A5FF",
      x"5FBB00BC",
      x"4BBE00BD",
      x"D58F40BF",
      x"B186705B",
      x"00BD00BC",
      x"40BF4BBE",
      x"7056D58A",
      x"00BCB186",
      x"4BBE00BD",
      x"D58540BF",
      x"B1867053",
      x"BC000003",
      x"000037C8",
      x"000037EC",
      x"000037FC",
      x"0000380A",
      x"40000000",
      x"0082B495",
      x"00000001",
      x"00000021",
      x"47311900",
      x"7D756A5A",
      x"6A757D7F",
      x"1931475A",
      x"B9CFE700",
      x"838B96A6",
      x"968B8381",
      x"E7CFB9A6",
      x"00001900",
      x"54BB00BC",
      x"55BE00BD",
      x"D58F40BF",
      x"B1867056",
      x"00BD00BC",
      x"40BF55BE",
      x"705BD58A",
      x"00BCB186",
      x"55BE00BD",
      x"D58540BF",
      x"B1867056",
      x"00BD00BC",
      x"40BF55BE",
      x"86705BD5",
      x"000000B1",
      x"B7000004",
      x"000037C8",
      x"00003860",
      x"00003870",
      x"0000387E",
      x"0000388C",
      x"4ABB00BC",
      x"78BE01BD",
      x"41E740BF",
      x"BCB19860",
      x"BE01BD00",
      x"E740BF78",
      x"B1987048",
      x"01BD00BC",
      x"40BF78BE",
      x"6C4CE782",
      x"00BCB198",
      x"78BE01BD",
      x"E78440BF",
      x"B1986C4F",
      x"01BD00BC",
      x"40BF78BE",
      x"6C53E786",
      x"00BCB198",
      x"78BE01BD",
      x"E78A40BF",
      x"B1986056",
      x"D0000006",
      x"000037C8",
      x"000038B4",
      x"000038C3",
      x"000038D0",
      x"000038DE",
      x"000038EC",
      x"000038FA",
      x"63BB00BC",
      x"5EBE00BD",
      x"D58F40BF",
      x"B1867864",
      x"00BD00BC",
      x"40BF5EBE",
      x"7862D58A",
      x"00BCB186",
      x"5EBE00BD",
      x"D58540BF",
      x"B1867860",
      x"00BD00BC",
      x"40BF5EBE",
      x"86505FD5",
      x"BD00BCB1",
      x"BF5EBE00",
      x"66D59440",
      x"BCB18678",
      x"BE00BD00",
      x"9840BF5E",
      x"7867DB81",
      x"0000B18C",
      x"B2000006",
      x"000037C8",
      x"00003928",
      x"00003938",
      x"00003946",
      x"00003954",
      x"00003961",
      x"0000396F",
      x"4ABB00BC",
      x"55BE02BD",
      x"D38440BF",
      x"B185786C",
      x"02BD00BC",
      x"40BF55BE",
      x"847060D3",
      x"000000B1",
      x"D0000002",
      x"000037C8",
      x"000039A0",
      x"000039B0",
      x"40000000",
      x"002F5658",
      x"00000000",
      x"00000520",
      x"3E483B0B",
      x"C6C3EB24",
      x"37350FDF",
      x"ADC0FF2A",
      x"321AE2BD",
      x"B0D61027",
      x"440DD9BD",
      x"D10D3346",
      x"32F4D1BE",
      x"053E5258",
      x"F6C9B5C4",
      x"1B3B4431",
      x"C9ACA5D4",
      x"23353503",
      x"C7AEB3F3",
      x"415134F1",
      x"C4BAE927",
      x"5C5115DF",
      x"B0DB264D",
      x"4619DDBB",
      x"B1F63045",
      x"26E5B8A2",
      x"CB0E2F3D",
      x"15D8B8A6",
      x"08374D4E",
      x"F8CFB7C6",
      x"3D58603A",
      x"CAAFBBFF",
      x"3E4E39FC",
      x"A9A0CE15",
      x"3C3C09CD",
      x"A9AEEC22",
      x"5639F6C7",
      x"B4E32244",
      x"561AE2BE",
      x"D61E4C64",
      x"1DE2B8AA",
      x"F02A4C4D",
      x"ECBA9DAF",
      x"06314529",
      x"DFB5A3C9",
      x"32535019",
      x"CFB1C501",
      x"5B663BFF",
      x"A9B7FA34",
      x"563A00CE",
      x"9DCE0C3C",
      x"400CD5A8",
      x"B0E71A41",
      x"38FECAA4",
      x"E217435B",
      x"1DE9BAB2",
      x"15466A57",
      x"EBBAA6D7",
      x"1F4F521C",
      x"C19AB2EE",
      x"2D4B28F2",
      x"B3A2CDFD",
      x"564F19E9",
      x"ACC8FD29",
      x"6A3805D3",
      x"B9F9275B",
      x"3902D7A7",
      x"D403345C",
      x"09DFAA9C",
      x"E70D4341",
      x"03D2A1B7",
      x"0C3E5C33",
      x"F3BAB3E7",
      x"3A6B541C",
      x"BFA5DB0E",
      x"4D5319F2",
      x"9AB7F113",
      x"4D24F5CA",
      x"A4D6F625",
      x"4B17F2B6",
      x"CDFB1D53",
      x"340ADAAB",
      x"FB1C5369",
      x"03E0ABBB",
      x"00295B37",
      x"E6B19FDB",
      x"033E3E06",
      x"DAA3BEEB",
      x"35582D05",
      x"BFB6EC06",
      x"66501AFA",
      x"AAE00B2F",
      x"5117F5C7",
      x"BDF50B44",
      x"20F5D2A0",
      x"DEF51B47",
      x"14F8BCAA",
      x"FD154B44",
      x"0BE1B1D4",
      x"1649622F",
      x"E4B4C3FC",
      x"20513302",
      x"BAA9E100",
      x"333704E9",
      x"ACC6F000",
      x"4C2705E0",
      x"BEF0052C",
      x"4919FDC7",
      x"E40A2858",
      x"15F5CFB6",
      x"F80A3847",
      x"F6D7ADC6",
      x"F914391B",
      x"F8C5B5E4",
      x"123D3911",
      x"E5BEDBFF",
      x"3D522C0A",
      x"C1CFFD15",
      x"412C02E4",
      x"B8E7021D",
      x"2A04E8C2",
      x"D1F50227",
      x"2004E1BA",
      x"F308253A",
      x"18FAD1CD",
      x"0927483C",
      x"F4D3C9EB",
      x"0E2E3514",
      x"D6BDD5FA",
      x"132612F6",
      x"CCC7EAFF",
      x"2F280FF5",
      x"CEE50016",
      x"3E2609E6",
      x"DFFE1736",
      x"2002E2CE",
      x"EE051F2F",
      x"01E6C7CD",
      x"F90B1C16",
      x"02DFCADF",
      x"0C242515",
      x"F7D9DEF7",
      x"28372B16",
      x"D5DBF50A",
      x"27210FF2",
      x"CBE5FD15",
      x"1405F5D3",
      x"DAF10417",
      x"1309F1D2",
      x"F1021B23",
      x"1B06E4DE",
      x"011A3229",
      x"00E0D9F1",
      x"09231F10",
      x"E3CCE0F8",
      x"131603FB",
      x"DDD8EFFE",
      x"241306FD",
      x"E0F0FE11",
      x"2B180FF3",
      x"EC000D2A",
      x"0F04EFD9",
      x"F7021A24",
      x"F7EFD2D8",
      x"FC0B1B06",
      x"FFEBD6EB",
      x"08201B01",
      x"00E5EBFE",
      x"1E2D180C",
      x"DFE3000A",
      x"251500F8",
      x"D0EF0310",
      x"13F4EEDE",
      x"E3FC061A",
      x"07F6F2DC",
      x"FC071823",
      x"0802EFE6",
      x"0B162A21",
      x"F7E8DDF7",
      x"0D202002",
      x"E3D2E102",
      x"151EFFE8",
      x"E3DDF607",
      x"2315F6ED",
      x"E7F30814",
      x"270EFEF4",
      x"EB071624",
      x"0EF5EADE",
      x"F80E1C26",
      x"EDDED5D7",
      x"05142110",
      x"E9E1DCEC",
      x"13222001",
      x"F1E9EE01",
      x"242A1800",
      x"DDE3FD13",
      x"291BFEE8",
      x"D2EB081C",
      x"1EFDDFD1",
      x"E4FC1123",
      x"10F0DBD6",
      x"FA0D2327",
      x"08F1E3E9",
      x"0A222F21",
      x"F0D9DBF4",
      x"162C270A",
      x"D0C7DFFE",
      x"232A0EEC",
      x"CCD9F408",
      x"301DFFE1",
      x"DDF5031D",
      x"2D11FBDF",
      x"E8011734",
      x"18FDDECE",
      x"F40A2A35",
      x"FCDCBFCD",
      x"FF19341F",
      x"F1CCC6EA",
      x"0E322E0B",
      x"E9D0E8FF",
      x"2C3E1D04",
      x"CAD4FB0A",
      x"3D2A08EE",
      x"B9E3001A",
      x"340CEFC7",
      x"D3F90930",
      x"1DFEDFB9",
      x"F804233F",
      x"0CF9D2D0",
      x"04184133",
      x"FDD8C0E8",
      x"0A334116",
      x"DEB2C6F8",
      x"1D4224FE",
      x"C4B6EA00",
      x"3D3809F2",
      x"C1E1000F",
      x"493B0BE5",
      x"B9E30319",
      x"4B1BFFD6",
      x"BEF70B39",
      x"2B00E0AC",
      x"E300204A",
      x"0DF2C0AB",
      x"FC10423F",
      x"00E1BBD7",
      x"09334F24",
      x"EFC0C6F5",
      x"1F4E390B",
      x"C4A8DA00",
      x"3C4615F6",
      x"AABFF30A",
      x"4D2900DC",
      x"BFE90029",
      x"4111F4C8",
      x"DBFD1A4A",
      x"2400D7BA",
      x"ED0A3B4E",
      x"08E2AEB9",
      x"FB224C33",
      x"F4C0A9D6",
      x"10424316",
      x"DDBBCEF1",
      x"354F2D05",
      x"C3C5E904",
      x"4E3F15EF",
      x"ABD1F820",
      x"4821FCC8",
      x"B8E4093D",
      x"3109DCAD",
      x"DAF92A4B",
      x"1DF4C7BF",
      x"F0194944",
      x"07D7C0D4",
      x"063C4E2F",
      x"E5B4BADF",
      x"244A3914",
      x"C1ADC8F0",
      x"404322F8",
      x"BFC9E00D",
      x"4C350EDB",
      x"CADBFC34",
      x"4322F2C9",
      x"C9EA204B",
      x"2D03CCB4",
      x"D3043C47",
      x"14DDB3B7",
      x"ED294636",
      x"F8C8C3CD",
      x"15454229",
      x"DCC9D1E0",
      x"3A4A3811",
      x"BDBFD2FE",
      x"463D21EC",
      x"B4BFE121",
      x"402C00C5",
      x"C7D0053E",
      x"3919DEC3",
      x"D1EF3047",
      x"2DFBD0D0",
      x"DC1A4743",
      x"0FD5BFC6",
      x"FA384435",
      x"E4BABAC5",
      x"2242381F",
      x"CDC6C6DE",
      x"40403101",
      x"D2D1D40A",
      x"473C1DE6",
      x"C5C9F133",
      x"3E2BF8C9",
      x"BBD21741",
      x"320ACEBA",
      x"C6F8363D",
      x"22E9C9C7",
      x"E3234039",
      x"07DED7CF",
      x"0C3C3E31",
      x"E6CECCD6",
      x"293A3318",
      x"CBC5C5ED",
      x"333121F2",
      x"D1CBD810",
      x"332B0BDE",
      x"DBD7FC2C",
      x"301EF8E1",
      x"D5EB1E35",
      x"2504E1D7",
      x"D7052C2F",
      x"0DE6D2CE",
      x"EF1C2A24",
      x"FADED7D4",
      x"0000000B",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000",
      x"00000000"
   );

begin

   process (clk) 
   begin
      if rising_edge(clk) then
         data <= rom(to_integer(unsigned(address)));
      end if;
   end process;

end architecture;
